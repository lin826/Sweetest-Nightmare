`ifndef _ROBOT_VH_
`define _ROBOT_VH_

`endif