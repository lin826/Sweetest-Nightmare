`ifndef _keyboard_vh_
`define _keyboard_vh_

`define ROW0 4'b1110
`define ROW1 4'b1101
`define ROW2 4'b1011
`define ROW3 4'b0111
	 
`define COL0 4'b0111
`define COL1 4'b1011
`define COL2 4'b1101
`define COL3 4'b1110

`define KEYCODE_EMPTY 16'hff

`define KEYCODE_F 16'b0111_1111_1111_1111
`define KEYCODE_E 16'b1011_1111_1111_1111
`define KEYCODE_D 16'b1101_1111_1111_1111
`define KEYCODE_C 16'b1110_1111_1111_1111

`define KEYCODE_B 16'b1111_0111_1111_1111
`define KEYCODE_3 16'b1111_1011_1111_1111
`define KEYCODE_6 16'b1111_1101_1111_1111
`define KEYCODE_9 16'b1111_1110_1111_1111

`define KEYCODE_A 16'b1111_1111_0111_1111
`define KEYCODE_2 16'b1111_1111_1011_1111
`define KEYCODE_5 16'b1111_1111_1101_1111
`define KEYCODE_8 16'b1111_1111_1110_1111

`define KEYCODE_0 16'b1111_1111_1111_0111
`define KEYCODE_1 16'b1111_1111_1111_1011
`define KEYCODE_4 16'b1111_1111_1111_1101
`define KEYCODE_7 16'b1111_1111_1111_1110

`endif

